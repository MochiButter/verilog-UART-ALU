module uart_echo
  (); 

endmodule
