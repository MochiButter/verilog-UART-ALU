`timescale 1ns / 1ps
module alu_state
  ();
  // controls the state of alu32.
endmodule
