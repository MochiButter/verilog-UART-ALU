`timescale 1ns/1ps
module top
  ();
  uart_echo #() ue_inst(

  );
endmodule 
